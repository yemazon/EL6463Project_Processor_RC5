----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:53:55 11/17/2017 
-- Design Name: 
-- Module Name:    instruction_memory - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;
--use STD.textio.all; -- Required for freading a file

entity instruction_memory is
	port (
		read_address: in STD_LOGIC_VECTOR (31 downto 0);
		instruction, last_instr_address: out STD_LOGIC_VECTOR (31 downto 0)
	);
end instruction_memory;

architecture Behavioral of instruction_memory is

	 type mem_array is array(0 to 157) of STD_LOGIC_VECTOR (31 downto 0);
    signal data_mem: mem_array := (
--		--|-Op-||Rs-||Rt-||------Im------|
--		--|----||---||---||--------------|
--	    "00000100000000110000000001001110",--ADDI 0 3 78
--
--		--|-Op-||Rs-||Rt-||------Im------|
--		--|----||---||---||--------------|
--		 "00000100000001000000000000011010",--ADDI 0 4 26
--
--		--|-Op-||Rs-||Rt-||------Im------|
--		--|----||---||---||--------------|
--		 "00000100000001010000000000000100",--ADDI 0 5 4
--        
--		-- OpCode|Rs ||Rt ||		imd		 |8
--	   -- |----||---||---||--------------|	
--		  "00011100000001100000000000000000", -- # lw
--		-- OpCode|Rs ||Rt ||		imd		 |8
--	   -- |----||---||---||--------------|	
--		  "00011100000001110000000000000001", -- # lw
--		  
--		--|-Op-||Rs-||Rt-||------Im------|1
--		--|----||---||---||--------------|
--		 "00000100000100010000000000000001",--ADDI 0 17 1
--
--		--|-Op-||Rs-||Rt-||------Im------|2
--		--|----||---||---||--------------|
--		 "00000100000100100000000000000010",--ADDI 0 18 2
--
--		--|-Op-||Rs-||Rt-||------Im------|3
--		--|----||---||---||--------------|
--		 "00000100000100110000000000000011",--ADDI 0 19 3
--		--|-Op-||Rs-||Rt-||------Im------|3
--		--|----||---||---||--------------|
--		 "00000100000101000000000000000100",--ADDI 0 20 4
--		-- Im 2
--		-- OpCode|Rs ||Rt ||		imd		 |4
--	   -- |----||---||---||--------------|
--        "00100001000001100000000000000000",
--		-- Im 3
--		-- OpCode|Rs ||Rt ||Rd ||Shm||Func|5
--	   -- |----||---||---||---||---||----|
--		  "00000000110001110011000000010000", -- # add
--		-- Im 3
--		-- OpCode|Rs ||Rt ||		imd		 |6
--	   -- |----||---||---||--------------|		  
--        "00000101000010000000000000000001", -- # andi
--		-- Im 4
--		-- OpCode|Rs ||Rt ||		imd		 |7
--	   -- |----||---||---||--------------|		  
--      --"00101101000001001111111111111100", -- # bne
--		  "00100101000001001111111111111100", -- # blt
--		-- Im 5
--		-- OpCode|Rs ||Rt ||		imd		 |8
--	   -- |----||---||---||--------------|	
--		  "00011100001011100000000000000000", -- # lw
--		-- Im 6
--		-- OpCode|Rs ||Rt ||Rd ||Shm||Func|9
--	   -- |----||---||---||---||---||----|
--		  "00000001011011000110100000010000", -- # add
--		-- Im 7
--		-- OpCode|Rs ||Rt ||Rd ||Shm||Func|10
--	   -- |----||---||---||---||---||----|
--		  "00000001101011100101100000010000", -- # add
--		-- Im 8
--		-- OpCode|Rs ||Rt ||		imd		 |11
--	   -- |----||---||---||--------------|	  
--		  "00010101011010110000000000000011",  -- # shl 3
--		-- Im 9
--		-- OpCode|Rs ||Rt ||		imd		 |12
--	   -- |----||---||---||--------------|
--		  "00100000001010110000000000000000",  -- # sw
--		-- Im 10
--		-- OpCode|Rs ||Rt ||		imd		 |13
--	   -- |----||---||---||--------------|	
--		  "00000100001000010000000000000001",  -- addi i++
--		-- Im 11
--		-- OpCode|Rs ||Rt ||		imd		 |14
--	   -- |----||---||---||--------------|	
--		  "00100100001001000000000000000010", -- blt
--		-- Im 12
--		-- OpCode|Rs ||Rt ||Rd ||Shm||Func|15
--	   -- |----||---||---||--------------| 
--		  "00001000001000010000000000011010", -- subi i-26
--		-- Im 13
--		-- OpCode|Rs ||Rt ||		imd		 |16
--	   -- |----||---||---||--------------|	
--		  "00101000000000001111111111111101", -- beq
--		-- Im 14
--		-- OpCode|Rs ||Rt ||		imd		 |17
--	   -- |----||---||---||--------------|	
--		  "00011100010011110000000000011010", -- lw
--		-- Im 15
--		-- OpCode|Rs ||Rt ||Rd ||Shm||Func|18
--	   -- |----||---||---||---||---||----|
--        "00000001011011000110100000010000", -- add A+B
--		-- Im 16
--		-- OpCode|Rs ||Rt ||Rd ||Shm||Func|19
--	   -- |----||---||---||---||---||----|
--        "00000001101011110110000000010000", -- add A + B + L[j]
--		-- Im 16.1
--		-- OpCode|Rs ||Rt ||		imd		 |20
--	   -- |----||---||---||--------------|	
--		  "00001101101011010000000000011111", -- andi
--		  
--		  
--		--|-Op-||Rs-||Rt-||------Im------|21
--		--|----||---||---||--------------|
--		 "00101000000011010000000000001100",--BEQ 0 13 12
--
--		--|-Op-||Rs-||Rt-||------Im------|22
--		--|----||---||---||--------------|
--		 "00100101101101000000000000000011",--BLT 13 20 3
--
--		--|-Op-||Rs-||Rt-||------Im------|23
--		--|----||---||---||--------------|
--		 "00001001101011010000000000000100",--SUBI 13 13 4
--
--		--|-Op-||Rs-||Rt-||------Im------|24
--		--|----||---||---||--------------|
--		 "00010101100011000000000000000100",--SHL 12 12 4
--
--		--|-Op-||Rs-||Rt-||------Im------|25
--		--|----||---||---||--------------|
--		 "00101000000000001111111111111011",--BEQ 0 0 -5
--
--		--|-Op-||Rs-||Rt-||------Im------|26
--		--|----||---||---||--------------|
--		  "00101110001011010000000000000010",--BNE 17 13 2
--
--		--|-Op-||Rs-||Rt-||------Im------|27
--		--|----||---||---||--------------|
--		 "00010101100011000000000000000001",--SHR 12 12 1
--
--		--|-Op-||Rs-||Rt-||------Im------|28
--		--|----||---||---||--------------|
--		  "00101000000000000000000000000101",--BEQ 0 0 5
--		--|-Op-||Rs-||Rt-||------Im------|29
--		--|----||---||---||--------------|
--		  "00101110010011010000000000000010",--BNE 18 13 2
--
--		--|-Op-||Rs-||Rt-||------Im------|30
--		--|----||---||---||--------------|
--		 "00010101100011000000000000000010",--SHR 12 12 2
--
--		--|-Op-||Rs-||Rt-||------Im------|
--		--|----||---||---||--------------|
--		  "00101000000000000000000000000010",--BEQ 0 0 2
--
--		--|-Op-||Rs-||Rt-||------Im------|
--		--|----||---||---||--------------|
--		  "00101110011011010000000000000001",--BNE 19 13 1
--
--		--|-Op-||Rs-||Rt-||------Im------|
--		--|----||---||---||--------------|
--		 "00010101100011000000000000000011",--SHR 12 12 3
--		-- Im 40
--		-- OpCode|Rs ||Rt ||		imd		 |
--	   -- |----||---||---||--------------|
--		  "00100000010011000000000000011010",  -- # sw
--		-- Im 41
--		-- OpCode|Rs ||Rt ||		imd		 |
--	   -- |----||---||---||--------------|	
--        "00000100010000100000000000000001",  -- # j++
--		-- Im 42
--		-- OpCode|Rs ||Rt ||		imd		 |
--	   -- |----||---||---||--------------|	
--		  "00100100010001010000000000000010", -- blt
--		-- Im 43
--		-- OpCode|Rs ||Rt ||Rd ||Shm||Func|
--	   -- |----||---||---||--------------| 
--		  "00001000010000100000000000000100", -- subi j-4
--		-- Im 44
--		-- OpCode|Rs ||Rt ||		imd		 |
--	   -- |----||---||---||--------------|	
--		  "00101000000000001111111111111101", -- beq
--      -- Im 45
--		-- OpCode|Rs ||Rt ||		imd		 |
--	   -- |----||---||---||--------------|	
--		  "00000110000100000000000000000001",  -- addi k++
--		-- Im 46
--		-- OpCode|Rs ||Rt ||		imd		 |
--	   -- |----||---||---||--------------|	
--		  "00100110000000111111111111011111", -- blt
--        "00000000000000000000000000000000",
--        "00000000000000000000000000000000", -- mem 30
--        "00000000000000000000000000000000", -- men 31
--		-- Im  
--		  "00000000000000000000000000000000", 
--        "00000000000000000000000000000000",
--		  "00000000000000000000000000000000",
--		  "00000000000000000000000000000000",
--        "00000000000000000000000000000000", 
--		  "00000000000000000000000000000000",
--        "00000000000000000000000000000000",
--		  "00000000000000000000000000000000",
--		  "00000000000000000000000000000000",
--        "00000000000000000000000000000000", 
--        "00000000000000000000000000000000",
--		  "00000000000000000000000000000000",
--        "00000000000000000000000000000000",
--        "00000000000000000000000000000000",
--		  "00000000000000000000000000000000"
    --|-Op-||Rs-||Rt-||------Im------|
    --|----||---||---||--------------|
      "00000100000000110000000001001110",--ADDI 0 3 78

    --|-Op-||Rs-||Rt-||------Im------|
    --|----||---||---||--------------|
     "00000100000001000000000000011010",--ADDI 0 4 26

    --|-Op-||Rs-||Rt-||------Im------|
    --|----||---||---||--------------|
     "00000100000001010000000000000100",--ADDI 0 5 4
        
    -- OpCode|Rs ||Rt ||    imd    |8
     -- |----||---||---||--------------|  
      "00011100000001100000000000000000", -- # lw
    -- OpCode|Rs ||Rt ||    imd    |8
     -- |----||---||---||--------------|  
      "00011100000001110000000000000001", -- # lw
      
    --|-Op-||Rs-||Rt-||------Im------|1
    --|----||---||---||--------------|
     "00000100000100010000000000000001",--ADDI 0 17 1

    --|-Op-||Rs-||Rt-||------Im------|2
    --|----||---||---||--------------|
     "00000100000100100000000000000010",--ADDI 0 18 2

    --|-Op-||Rs-||Rt-||------Im------|3
    --|----||---||---||--------------|
     "00000100000100110000000000000011",--ADDI 0 19 3
    --|-Op-||Rs-||Rt-||------Im------|3
    --|----||---||---||--------------|
     "00000100000101000000000000000100",--ADDI 0 20 4
    -- Im 2
    -- OpCode|Rs ||Rt ||    imd    |4
     -- |----||---||---||--------------|
        "00100001000001100000000000000000",
    -- Im 3
    -- OpCode|Rs ||Rt ||Rd ||Shm||Func|5
     -- |----||---||---||---||---||----|
      "00000000110001110011000000010000", -- # add
    -- Im 3
    -- OpCode|Rs ||Rt ||    imd    |6
     -- |----||---||---||--------------|      
        "00000101000010000000000000000001", -- # andi
    -- Im 4
    -- OpCode|Rs ||Rt ||    imd    |7
     -- |----||---||---||--------------|      
      --"00101101000001001111111111111100", -- # bne
      "00100101000001001111111111111100", -- # blt
    -- Im 5
    -- OpCode|Rs ||Rt ||    imd    |8
     -- |----||---||---||--------------|  
      "00011100001011100000000000000000", -- # lw
    -- Im 6
    -- OpCode|Rs ||Rt ||Rd ||Shm||Func|9
     -- |----||---||---||---||---||----|
      "00000001011011000110100000010000", -- # add
    -- Im 7
    -- OpCode|Rs ||Rt ||Rd ||Shm||Func|10
     -- |----||---||---||---||---||----|
      "00000001101011100101100000010000", -- # add
    -- Im 8
    -- OpCode|Rs ||Rt ||    imd    |11
     -- |----||---||---||--------------|    
      "00010101011010110000000000000011",  -- # shl 3
    -- Im 9
    -- OpCode|Rs ||Rt ||    imd    |12
     -- |----||---||---||--------------|
      "00100000001010110000000000000000",  -- # sw
    -- Im 10
    -- OpCode|Rs ||Rt ||    imd    |13
     -- |----||---||---||--------------|  
      "00000100001000010000000000000001",  -- addi i++
    -- Im 11
    -- OpCode|Rs ||Rt ||    imd    |14
     -- |----||---||---||--------------|  
      "00100100001001000000000000000010", -- blt
    -- Im 12
    -- OpCode|Rs ||Rt ||Rd ||Shm||Func|15
     -- |----||---||---||--------------| 
      "00001000001000010000000000011010", -- subi i-26
    -- Im 13
    -- OpCode|Rs ||Rt ||    imd    |16
     -- |----||---||---||--------------|  
      "00101000000000001111111111111101", -- beq
    -- Im 14
    -- OpCode|Rs ||Rt ||    imd    |17
     -- |----||---||---||--------------|  
      "00011100010011110000000000011010", -- lw
    -- Im 15
    -- OpCode|Rs ||Rt ||Rd ||Shm||Func|18
     -- |----||---||---||---||---||----|
        "00000001011011000110100000010000", -- add A+B
    -- Im 16
    -- OpCode|Rs ||Rt ||Rd ||Shm||Func|19
     -- |----||---||---||---||---||----|
        "00000001101011110110000000010000", -- add A + B + L[j]
    -- Im 16.1
    -- OpCode|Rs ||Rt ||    imd    |20
     -- |----||---||---||--------------|  
      "00001101101011010000000000011111", -- andi
      
      
    --|-Op-||Rs-||Rt-||------Im------|21
    --|----||---||---||--------------|
     "00101000000011010000000000001100",--BEQ 0 13 12

    --|-Op-||Rs-||Rt-||------Im------|22
    --|----||---||---||--------------|
     "00100101101101000000000000000011",--BLT 13 20 3

    --|-Op-||Rs-||Rt-||------Im------|23
    --|----||---||---||--------------|
     "00001001101011010000000000000100",--SUBI 13 13 4

    --|-Op-||Rs-||Rt-||------Im------|24
    --|----||---||---||--------------|
     "00010101100011000000000000000100",--SHL 12 12 4

    --|-Op-||Rs-||Rt-||------Im------|25
    --|----||---||---||--------------|
     "00101000000000001111111111111011",--BEQ 0 0 -5

    --|-Op-||Rs-||Rt-||------Im------|26
    --|----||---||---||--------------|
      "00101110001011010000000000000010",--BNE 17 13 2

    --|-Op-||Rs-||Rt-||------Im------|27
    --|----||---||---||--------------|
     "00010101100011000000000000000001",--SHR 12 12 1

    --|-Op-||Rs-||Rt-||------Im------|28
    --|----||---||---||--------------|
      "00101000000000000000000000000101",--BEQ 0 0 5
    --|-Op-||Rs-||Rt-||------Im------|29
    --|----||---||---||--------------|
      "00101110010011010000000000000010",--BNE 18 13 2

    --|-Op-||Rs-||Rt-||------Im------|30
    --|----||---||---||--------------|
     "00010101100011000000000000000010",--SHR 12 12 2

    --|-Op-||Rs-||Rt-||------Im------|
    --|----||---||---||--------------|
      "00101000000000000000000000000010",--BEQ 0 0 2

    --|-Op-||Rs-||Rt-||------Im------|
    --|----||---||---||--------------|
      "00101110011011010000000000000001",--BNE 19 13 1

    --|-Op-||Rs-||Rt-||------Im------|
    --|----||---||---||--------------|
     "00010101100011000000000000000011",--SHR 12 12 3
    -- Im 40
    -- OpCode|Rs ||Rt ||    imd    |
     -- |----||---||---||--------------|
      "00100000010011000000000000011010",  -- # sw
    -- Im 41
    -- OpCode|Rs ||Rt ||    imd    |
     -- |----||---||---||--------------|  
        "00000100010000100000000000000001",  -- # j++
    -- Im 42
    -- OpCode|Rs ||Rt ||    imd    |
     -- |----||---||---||--------------|  
      "00100100010001010000000000000010", -- blt
    -- Im 43
    -- OpCode|Rs ||Rt ||Rd ||Shm||Func|
     -- |----||---||---||--------------| 
      "00001000010000100000000000000100", -- subi j-4
    -- Im 44
    -- OpCode|Rs ||Rt ||    imd    |
     -- |----||---||---||--------------|  
      "00101000000000001111111111111101", -- beq
      -- Im 45
    -- OpCode|Rs ||Rt ||    imd    |
     -- |----||---||---||--------------|  
      "00000110000100000000000000000001",  -- addi k++
    -- Im 46
    -- OpCode|Rs ||Rt ||    imd    |
     -- |----||---||---||--------------|  
      "00100110000000111111111111011111", -- blt
		  
		  
		  
		  		----encrypt

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00011100000000010000000000011110",--LW 0 1 30

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00011100000000100000000000011111",--LW 0 2 31

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00011100000010010000000000000000",--LW 0 9 0

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00000100000010110000000000000001",--ADDI 0 11 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00000100000011000000000000000010",--ADDI 0 12 2

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00000100000011010000000000000011",--ADDI 0 13 3

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000001010010000100000010000",--ADD 1 9 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00011100000010010000000000000001",--LW 0 9 1

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000010010010001000000010000",--ADD 2 9 2

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00000100000000110000000000000010",--ADDI 0 3 2

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00000100000010000000000000011010",--ADDI 0 8 26

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000001000010010000000010100",--NOR 1 1 4

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000010000100010100000010100",--NOR 2 2 5

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000001001010011000000010010",--AND 1 5 6

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000010001000011100000010010",--AND 2 4 7

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000110001110000100000010011",--OR 6 7 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00001100010010100000000000011111",--ANDI 2 10 31

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00101001010000000000000000001010",--BEQ 10 0 10

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00101001010010110000000000001000",--BEQ 10 11 8

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00101001010011000000000000000110",--BEQ 10 12 6

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00101001010011010000000000000100",--BEQ 10 13 4

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00010100001000010000000000000100",--SHL 1 1 4

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00001001010010100000000000000100",--SUBI 10 10 4

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00101101010000001111111111111010",--BNE 10 0 -6
  
--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00101001010000000000000000000011",--BEQ 10 0 3

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00010100001000010000000000000001",--SHL 1 1 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00010100001000010000000000000001",--SHL 1 1 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00010100001000010000000000000001",--SHL 1 1 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00011100011010010000000000000000",--LW 3 9 0

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000001010010000100000010000",--ADD 1 9 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00000100011000110000000000000001",--ADDI 3 3 1

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000001000010010000000010100",--NOR 1 1 4

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000010000100010100000010100",--NOR 2 2 5

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000001001010011000000010010",--AND 1 5 6

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000010001000011100000010010",--AND 2 4 7

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000110001110001000000010011",--OR 6 7 2

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00001100001010100000000000011111",--ANDI 1 10 31

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00101001010000000000000000001010",--BEQ 10 0 10

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00101001010010110000000000001000",--BEQ 10 11 8

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00101001010011000000000000000110",--BEQ 10 12 6

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00101001010011010000000000000100",--BEQ 10 13 4

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00010100010000100000000000000100",--SHL 2 2 4

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00001001010010100000000000000100",--SUBI 10 10 4

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00101101010000001111111111111010",--BNE 10 0 -6
  
--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00101001010000000000000000000011",--BEQ 10 0 3
  

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00010100010000100000000000000001",--SHL 2 2  1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00010100010000100000000000000001",--SHL 2 2 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00010100010000100000000000000001",--SHL 2 2 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00011100011010010000000000000000",--LW 3 9 0

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
  "00000000010010010001000000010000",--ADD 2 9 2

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00000100011000110000000000000001",--ADDI 3 3 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101100011010001111111111010111",--BNE 3 8 -41

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
  "00100000000000010000000000100000",--SW 0 1 32

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------| --SW 0 2 33
  "00100000000000100000000000100001",
  
  -----decrypt
  --|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011100000000010000000000011110",--LW 0 1 30

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011100000000100000000000011111",--LW 0 2 31

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00000100000000110000000000011001",--ADDI 0 3 25

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00000100000010100000000000000001",--ADDI 0 10 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00000100000010110000000000000100",--ADDI 0 11 4

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00000100000011000000000000000011",--ADDI 0 12 3

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00000100000011010000000000000010",--ADDI 0 13 2

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00000100000011100000000000000001",--ADDI 0 14 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011100011010000000000000000000",--LW 3 8 0

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000010010000001000000010001",--SUB 2 8 2 

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00001100001010010000000000011111",--ANDI 1 9 31

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101001001000000000000000001010",--BEQ 9 0 10
----------------------------------------------------------
--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101001100010010000000000000110",--BEQ 12 9 6

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101001101010010000000000000110",--BEQ 13 9 6

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101001110010010000000000000110",--BEQ 14 9 6

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011000010000100000000000000100",--SHR 2 2 4

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00001001001010010000000000000100",--SUBI 9 9 4

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101100000010011111111111111010",--BNE 0 9 -6

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101000000010010000000000000011",--BEQ 0 9 3

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011000010000100000000000000001",--SHR 2 2 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011000010000100000000000000001",--SHR 2 2 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011000010000100000000000000001",--SHR 2 2 1

----------------------------------------------------------
--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000001000010010000000010100",--NOR 1 1 4

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000010000100010100000010100",--NOR 2 2 5

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000001001010011000000010010",--AND 1 5 6

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000010001000011100000010010",--AND 2 4 7

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000110001110001000000010011",--OR 6 7 2

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00001000011000110000000000000001",--SUBI 3 3 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011100011010000000000000000000",--LW 3 8 0

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000001010000000100000010001",--SUB 1 8 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00001100010010010000000000011111",--ANDI 2 9 31

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101001001000000000000000001010",--BEQ 9 0 10
----------------------------------------------------------
--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101001100010010000000000000110",--BEQ 12 9 6

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101001101010010000000000000110",--BEQ 13 9 6

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101001110010010000000000000110",--BEQ 14 9 6

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011000001000010000000000000100",--SHR 1 1 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00001001001010010000000000000100",--SUBI 9 9 4

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101100000010011111111111111010",--BNE 0 9 -6

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101000000010010000000000000011",--BEQ 0 9 3

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011000001000010000000000000001",--SHR 1 1 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011000001000010000000000000001",--SHR 1 1 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011000001000010000000000000001",--SHR 1 1 1
----------------------------------------------------------
--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000001000010010000000010100",--NOR 1 1 4

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000010000100010100000010100",--NOR 2 2 5

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000001001010011000000010010",--AND 1 5 6

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000010001000011100000010010",--AND 2 4 7

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000110001110000100000010011",--OR 6 7 2

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00001000011000110000000000000001",--SUBI 3 3 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00101100011010101111111111010111",--BNE 3 10 -41

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011100011010000000000000000000",--LW 3 8 0

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-|
--|----||---||---||---||---||----|
 "00000000010010000001000000010001",--SUB 2 8 2

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00001000011000110000000000000001",--SUBI 3 3 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00011100011010000000000000000000",--LW 3 8 0

--|-Op-||Rs-||Rt-||Rd-||Sh-||-Fc-| 
--|----||---||---||---||---||----|
 "00000000001010000000100000010001",--SUB 1 8 1

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00100000000000010000000000100010",--SW 0 1 34

--|-Op-||Rs-||Rt-||------Im------|
--|----||---||---||--------------|
 "00100000000000100000000000100011",
 "00101000000000001111111111111111", -- beq
  "00000000000000000000000000000000"
    );

begin

    instruction <= data_mem(to_integer(unsigned(read_address(31 downto 2))));

end Behavioral;

